module font_rom ( input [10:0]	addr,
						//output [15:0]	data
						output [23:0] data
					 );

	parameter ADDR_WIDTH = 11;
   //parameter DATA_WIDTH =  16;
	parameter DATA_WIDTH = 24;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
//	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
parameter [0:285][DATA_WIDTH-1:0] ROM = {
		  
		  24'b000000000000000000000000, // 0
        24'b000000000000000000000000, // 1
        24'b000000000000000000000000, // 2
        24'b000000000000000000000000, // 3
        24'b000000000000000000000000, // 4
        24'b000000000000000000000000, // 5
        24'b000000000000000000000000, // 6
        24'b000000000000000000000000, // 7
        24'b000000000000000000000000, // 8
        24'b000000000000000000000000, // 9
        24'b000000000000000000000000, // 10
        24'b000000000000000000000000, // 11
        24'b000000000000000000000000, // 12
        24'b000000000000000000000000, // 13
        24'b000000000000000000000000, // 14
        24'b000000000000000000000000, // 15
        24'b000000000000000000000000, // 16
        24'b000000000000000000000000, // 17
        24'b000000000000000000000000, // 18
        24'b000000000000000000000000, // 19
        24'b000000000000000000000000, // 20
        24'b000000000000000000000000, // 21
		  
		  // code x01 (facing upwards)
		  //  010101010101010101010101
		  24'b000000000000000000000000, // 0
        24'b001110000000000000011110, // 1
        24'b111110001111111100011111, // 2
        24'b111110110111111011011111, // 3
        24'b011110100111111001011110, // 4
        24'b011110111111111111011110, // 5
        24'b011111111111111111111110, // 6
        24'b011111111111111111111110, // 7
        24'b001111111111111111111100, // 8
        24'b000001111111111111100000, // 9
		  24'b000001111111111111100000, // 10
		  24'b000001111111111111100000, // 11
		  24'b000001111111111111100000, // 12
		  24'b000001111111111111100000, // 13
		  24'b001111111111111111111100, // 14
        24'b011111111111111111111110, // 15
        24'b011111111111111111111110, // 16
        24'b011111111111111111111110, // 17
        24'b111110111111111111011111, // 18
        24'b111110001111111100011111, // 19
        24'b011110000000000000011110, // 20
        24'b000000000000000000000000, // 21
		  
		  // code x02 (facing downwards)
		  //  010101010101010101010101
		  24'b000000000000000000000000, // 0
		  24'b011110000111111000011110, // 1
		  24'b111110001111111100011111, // 2
		  24'b111110111111111111011111, // 3
		  24'b011111111111111111111110, // 4
		  24'b011111111111111111111110, // 5
		  24'b011111111111111111111110, // 6
		  24'b001111111111111111111100, // 7
		  24'b000001111111111111100000, // 8
		  24'b000001111111111111100000, // 9
		  24'b000001111111111111100000, // 10
		  24'b000001111111111111100000, // 11
		  24'b000001111111111111100000, // 12 
		  24'b001111111111111111111100, // 13 
		  24'b011111111111111111111110, // 14
		  24'b011111111111111111111110, // 15
		  24'b011110111111111111011110, // 16
		  24'b011110100111111001011110, // 17
		  24'b111110110111111011011111, // 18
		  24'b111110001111111100011111, // 19
		  24'b011110000000000000011110, // 20
		  24'b000000000000000000000000, // 21
		  
		  
		  // code x03 (facing right for some reason even though it's coded to look left)
		  //  010101010101010101010101
		  24'b011111110000000001111110, // 0
		  24'b111111111000000011111111, // 1
		  24'b111111111000000011111111, // 2
		  24'b111111111000000011111111, // 3
		  24'b000000111111111111110000, // 4
		  24'b000111111111111111111000, // 5
		  24'b000101111111111111111000, // 6
		  24'b001001111111111111111100, // 7
		  24'b001111111111111111111110, // 8
		  24'b001111111111111111111110, // 9
		  24'b001111111111111111111110, // 10
		  24'b001111111111111111111110, // 11
		  24'b001111111111111111111110, // 12
		  24'b001111111111111111111110, // 13
		  24'b001001111111111111111100, // 14
		  24'b000101111111111111111000, // 15
		  24'b000111111111111111111000, // 16
		  24'b000000111111111111110000, // 17
		  24'b111111111000000011111111, // 18
		  24'b111111111000000011111111, // 19
		  24'b111111111000000011111111, // 20
		  24'b011111110000000001111110, // 21
		  
		  // code x04 (facing left for some reason even though it's coded to look right)
		  //  010101010101010101010101
		  24'b011111100000000011111110, // 0
		  24'b111111110000000111111111, // 1
		  24'b111111110000000111111111, // 2
		  24'b111111110000000111111111, // 3
		  24'b000011111111111111000000, // 4
		  24'b000111111111111111111000, // 5
		  24'b000111111111111111101000, // 6
		  24'b001111111111111111100100, // 7
		  24'b011111111111111111111100, // 8
		  24'b011111111111111111111100, // 9
		  24'b011111111111111111111100, // 10
		  24'b011111111111111111111100, // 11
		  24'b011111111111111111111100, // 12
		  24'b011111111111111111111100, // 13
		  24'b001111111111111111100100, // 14
		  24'b000111111111111111101000, // 15
		  24'b000111111111111111111000, // 16
		  24'b000011111111111111000000, // 17
		  24'b111111110000000111111111, // 18
		  24'b111111110000000111111111, // 19
		  24'b111111110000000111111111, // 20
		  24'b011111100000000011111110, // 21
		  
		  // code x05
		  24'b000000000000000000000000, // 0			
        24'b000000000000000000000000, // 1
        24'b000000000000000000000000, // 2		  
        24'b000000000000000000000000, // 3
        24'b000000000000000000000000, // 4
        24'b000000000111110000000000, // 5	  *****
        24'b000000001100011000000000, // 6	 **   **
        24'b000000001100011000000000, // 7 	**   **
        24'b000000000110000000000000, // 8	  **
        24'b000000000011100000000000, // 9	   ***
        24'b000000000000110000000000, // 10	     **
        24'b000000000000011000000000, // 11	      **
        24'b000000001100011000000000, // 12	 **   **
        24'b000000001100011000000000, // 13	 **   **
        24'b000000000111110000000000, // 14	  *****
        24'b000000000000000000000000, // 15
        24'b000000000000000000000000, // 16
        24'b000000000000000000000000, // 17
        24'b000000000000000000000000, // 18
		  24'b000000000000000000000000, // 19
        24'b000000000000000000000000, // 20	  
		  24'b000000000000000000000000, // 21	

         // code x06		
        24'b000000000000000000000000, // 0
        24'b000000000000000000000000, // 1
        24'b000000000000000000000000, // 2		  
        24'b000000000000000000000000, // 3
        24'b000000000000000000000000, // 4
        24'b000000000011110000000000, // 5	   ****
        24'b000000000110011000000000, // 6	  **  **
        24'b000000001100001000000000, // 7	 **    *
        24'b000000001100000000000000, // 8	 **
        24'b000000001100000000000000, // 9	 **
        24'b000000001100000000000000, // 10	 **
        24'b000000001100000000000000, // 11	 **
        24'b000000001100001000000000, // 12	 **    *
        24'b000000000110011000000000, // 13	  **  **
        24'b000000000011110000000000, // 14	   ****
        24'b000000000000000000000000, // 15
        24'b000000000000000000000000, // 16
        24'b000000000000000000000000, // 17
        24'b000000000000000000000000, // 18
		  24'b000000000000000000000000, // 19
		  24'b000000000000000000000000, // 20
		  24'b000000000000000000000000, // 21


         // code x07			
        24'b000000000000000000000000, // 0
        24'b000000000000000000000000, // 1
        24'b000000000000000000000000, // 2		  
        24'b000000000000000000000000, // 3
        24'b000000000000000000000000, // 4
        24'b000000000111110000000000, // 5	  *****
        24'b000000001100011000000000, // 6	 **   **
        24'b000000001100011000000000, // 7	 **   **
        24'b000000001100011000000000, // 8	 **   **
        24'b000000001100011000000000, // 9	 **   **
        24'b000000001100011000000000, // 10	 **   **
        24'b000000001100011000000000, // 11	 **   **
        24'b000000001100011000000000, // 12	 **   **
        24'b000000001100011000000000, // 13	 **   **
        24'b000000000111110000000000, // 14	  *****
        24'b000000000000000000000000, // 15
        24'b000000000000000000000000, // 16
        24'b000000000000000000000000, // 17
        24'b000000000000000000000000, // 18
        24'b000000000000000000000000, // 19
		  24'b000000000000000000000000, // 20
        24'b000000000000000000000000, // 21
		  

         // code x08
        24'b000000000000000000000000, // 0
        24'b000000000000000000000000, // 1
        24'b000000000000000000000000, // 2		  
        24'b000000000000000000000000, // 3
        24'b000000000000000000000000, // 4
        24'b000000001111110000000000, // 5	 ******
        24'b000000000110011000000000, // 6	  **  **
        24'b000000000110011000000000, // 7	  **  **
        24'b000000000110011000000000, // 8	  **  **
        24'b000000000111110000000000, // 9	  *****
        24'b000000000110110000000000, // 10	  ** **
        24'b000000000110011000000000, // 11	  **  **
        24'b000000000110011000000000, // 12	  **  **
        24'b000000000110011000000000, // 13	  **  **
        24'b000000001110011000000000, // 14	 ***  **
        24'b000000000000000000000000, // 15
        24'b000000000000000000000000, // 16
        24'b000000000000000000000000, // 17
        24'b000000000000000000000000, // 18
        24'b000000000000000000000000, // 19
		  24'b000000000000000000000000, // 20
        24'b000000000000000000000000, // 21
	

         // code x09
        24'b000000000000000000000000, // 0
        24'b000000000000000000000000, // 1
        24'b000000000000000000000000, // 2		  
        24'b000000000000000000000000, // 3
        24'b000000000000000000000000, // 4
        24'b000000001111111000000000, // 5	 *******
        24'b000000000110011000000000, // 6	  **  **
        24'b000000000110001000000000, // 7	  **   *
        24'b000000000110100000000000, // 8	  ** *
        24'b000000000111100000000000, // 9	  ****
        24'b000000000110100000000000, // 10	  ** *
        24'b000000000110000000000000, // 11	  **
        24'b000000000110001000000000, // 12	  **   *
        24'b000000000110011000000000, // 13	  **  **
        24'b000000001111111000000000, // 14	 *******
        24'b000000000000000000000000, // 15
        24'b000000000000000000000000, // 16
        24'b000000000000000000000000, // 17
        24'b000000000000000000000000, // 18
        24'b000000000000000000000000, // 19
		  24'b000000000000000000000000, // 20
        24'b000000000000000000000000, // 21
	

         // code x0a		  
        24'b000000000000000000000000, // 0
        24'b000000000000000000000000, // 1
        24'b000000000000000000000000, // 2		  
        24'b000000000000000000000000, // 3
        24'b000000000000000000000000, // 4
        24'b000000000000000000000000, // 5
        24'b000000000000000000000000, // 6
        24'b000000000001100000000000, // 7	    **
        24'b000000000001100000000000, // 8	    **
        24'b000000000000000000000000, // 9
        24'b000000000000000000000000, // 10
        24'b000000000000000000000000, // 11
        24'b000000000001100000000000, // 12	    **
        24'b000000000001100000000000, // 13	    **
        24'b000000000000000000000000, // 14
        24'b000000000000000000000000, // 15
        24'b000000000000000000000000, // 16
        24'b000000000000000000000000, // 17
        24'b000000000000000000000000, // 18
        24'b000000000000000000000000, // 19
		  24'b000000000000000000000000, // 20
        24'b000000000000000000000000, // 21
		
        
		  // code x0b
        24'b000000000000000000000000, // 0
        24'b000000000000000000000000, // 1
        24'b000000000000000000000000, // 2		  
        24'b000000000000000000000000, // 3
        24'b000000000000000000000000, // 4
        24'b000000000111110000000000, // 5	  *****
        24'b000000001100011000000000, // 6	 **   **
        24'b000000001100011000000000, // 7	 **   **
        24'b000000001100111000000000, // 8	 **  ***
        24'b000000001101111000000000, // 9	 ** ****
        24'b000000001111011000000000, // 10	 **** **
        24'b000000001110011000000000, // 11	 ***  **
        24'b000000001100011000000000, // 12	 **   **
        24'b000000001100011000000000, // 13	 **   **
        24'b000000000111110000000000, // 14	  *****
        24'b000000000000000000000000, // 15
        24'b000000000000000000000000, // 16
        24'b000000000000000000000000, // 17
        24'b000000000000000000000000, // 18
        24'b000000000000000000000000, // 19
		  24'b000000000000000000000000, // 20
        24'b000000000000000000000000, // 21
		  
		  // code x0c
		  24'b111111111111111111111111, // 0
		  24'b111111111111111111111111, // 1
		  24'b111111111111111111111111, // 2
		  24'b111111111111111111111111, // 3
		  24'b111111111111111111111111, // 4
		  24'b111111111111111111111111, // 5
		  24'b111111111111111111111111, // 6
		  24'b111111111111111111111111, // 7
		  24'b111111111111111111111111, // 8
		  24'b111111111111111111111111, // 9
		  24'b111111111111111111111111, // 10
		  24'b111111111111111111111111, // 11
		  24'b111111111111111111111111, // 12
		  24'b111111111111111111111111, // 13
		  24'b111111111111111111111111, // 14
		  24'b111111111111111111111111, // 15
		  24'b111111111111111111111111, // 16
		  24'b111111111111111111111111, // 17
		  24'b111111111111111111111111, // 18
		  24'b111111111111111111111111, // 19
		  24'b111111111111111111111111, // 20
		  24'b111111111111111111111111 // 21 
		  
        };		  

	assign data = ROM[addr];

endmodule  